////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : apb_seq_pkg
// Description    : Dummy seq_pkg which can be used to create new seq_pkg
///////////////////////////////////////////////////////////////////////
package apb_seq_pkg;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	`include "apb_mst_seq_item.sv"
	`include "apb_slv_seq_item.sv"
	`include "apb_mst_seq_lib.sv"
	`include "apb_slv_seq_lib.sv"
endpackage