////////////////////////////////////////////////////////////////////////
// Developer Name : Mohsan Naeem 
// Contact info   : mohsannaeem1576@gmail.com
// Module Name    : apb_env_pkg
// Description    : Dummy env_pkg which can be used to create new env_pkg
///////////////////////////////////////////////////////////////////////
package apb_env_pkg;
   import uvm_pkg::*;
   `include "uvm_macros.svh"
   import apb_seq_pkg::*;
   `include "apb_agent_config.sv"
   `include "apb_env_config.sv"
   `include "apb_mst_sequencer.sv"
   `include "apb_mst_driver.sv"
   `include "apb_mst_monitor.sv"
   `include "apb_mst_agent.sv"
   `include "apb_slv_sequencer.sv"
   `include "apb_slv_driver.sv"
   `include "apb_slv_monitor.sv"
   `include "apb_slv_agent.sv"
   `include "apb_env.sv"
endpackage